module 7-segment
(
input clk,
input button,

output led1;
output led2;
output led3;
output led4;
output led5;
output led6;
output led7;
output led8;

output control_led1;
output control_led2;
output control_led3;
output control_led4;
);