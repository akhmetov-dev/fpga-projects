// unsaved_tb.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module unsaved_tb (
	);

	wire    unsaved_inst_clk_bfm_clk_clk;       // unsaved_inst_clk_bfm:clk -> [unsaved_inst:clk_clk, unsaved_inst_reset_bfm:clk]
	wire    unsaved_inst_reset_bfm_reset_reset; // unsaved_inst_reset_bfm:reset -> unsaved_inst:reset_reset_n

	unsaved unsaved_inst (
		.clk_clk       (unsaved_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (unsaved_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) unsaved_inst_clk_bfm (
		.clk (unsaved_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) unsaved_inst_reset_bfm (
		.reset (unsaved_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (unsaved_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
